package shared_pkg;

  bit    test_finished = 0;
  int    error_count = 0;
  int    correct_count = 0;
  event  sample_event;

endpackage
